module controlpath();
loduuu
endmodule