module Instruction_Memory(
    input [31:0] address,
    output [31:0] data
);
    reg [31:0] RAM [0:96];
    assign data = RAM[address[7:2]];
    initial begin
        /*mem[0] = 32'h000000B3;  
        mem[1] = 32'h00000233;  
        mem[2] = 32'h00A08113;  
        mem[3] = 32'h000081B3;  
        mem[4] = 32'h00218863;  
        mem[5] = 32'h00418233;  
        //mem[6] = 32'hFE21CCE3;
        mem[6] = 32'h00118193;
        mem[7] = 32'hfe000ae3; 
        mem[8] = 32'h000200b3;*/
        RAM[0] = 32'h00000093; // addi x1, x0, 0
    RAM[1] = 32'h00100113; // addi x2, x0, 1

    // Store first two numbers to memory 0(x0) and 4(x0)
    RAM[2] = 32'h00102023; // sw x1, 0(x0) = 0
    RAM[3] = 32'h00202223; // sw x2, 4(x0) = 1

    // Generate Fibonacci numbers (fully unrolled, storing each result to memory)
    RAM[4]  = 32'h002081B3; // add x3, x1, x2 => 0+1=1
    RAM[5]  = 32'h00302423; // sw x3, 8(x0) => 1
    RAM[6]  = 32'h002000B3; // add x1, x0, x2 => x1=1
    RAM[7]  = 32'h00300133; // add x2, x0, x3 => x2=1

    RAM[8]  = 32'h002081B3; // add x3, x1, x2 => 1+1=2
    RAM[9]  = 32'h00302623; // sw x3, 12(x0) => 2
    RAM[10] = 32'h002000B3; // add x1, x0, x2 => x1=1
    RAM[11] = 32'h00300133; // add x2, x0, x3 => x2=2

    RAM[12] = 32'h002081B3; // add x3, x1, x2 => 1+2=3
    RAM[13] = 32'h00302823; // sw x3, 16(x0) => 3
    RAM[14] = 32'h002000B3; // add x1, x0, x2 => x1=2
    RAM[15] = 32'h00300133; // add x2, x0, x3 => x2=3

    RAM[16] = 32'h002081B3; // add x3, x1, x2 => 2+3=5
    RAM[17] = 32'h00302A23; // sw x3, 20(x0) => 5
    RAM[18] = 32'h002000B3; // add x1, x0, x2 => x1=3
    RAM[19] = 32'h00300133; // add x2, x0, x3 => x2=5

    RAM[20] = 32'h002081B3; // add x3, x1, x2 => 3+5=8
    RAM[21] = 32'h00302C23; // sw x3, 24(x0) => 8
    RAM[22] = 32'h002000B3; // add x1, x0, x2 => x1=5
    RAM[23] = 32'h00300133; // add x2, x0, x3 => x2=8

    RAM[24] = 32'h002081B3; // add x3, x1, x2 => 5+8=13
    RAM[25] = 32'h00302E23; // sw x3, 28(x0) => 13
    RAM[26] = 32'h002000B3; // add x1, x0, x2 => x1=8
    RAM[27] = 32'h00300133; // add x2, x0, x3 => x2=13

    RAM[28] = 32'h002081B3; // add x3, x1, x2 => 8+13=21
    RAM[29] = 32'h003020A3; // sw x3, 32(x0) => 21
    RAM[30] = 32'h002000B3; // add x1, x0, x2 => x1=13
    RAM[31] = 32'h00300133; // add x2, x0, x3 => x2=21

    RAM[32] = 32'h002081B3; // add x3, x1, x2 => 13+21=34
    RAM[33] = 32'h003022A3; // sw x3, 36(x0) => 34
    RAM[34] = 32'h002000B3; // add x1, x0, x2 => x1=21
    RAM[35] = 32'h00300133; // add x2, x0, x3 => x2=34

    RAM[36] = 32'h002081B3; // add x3, x1, x2 => 21+34=55
    RAM[37] = 32'h003024A3; // sw x3, 40(x0) => 55
    RAM[38] = 32'h002000B3; // add x1, x0, x2 => x1=34
    RAM[39] = 32'h00300133; // add x2, x0, x3 => x2=55

    RAM[40] = 32'h002081B3; // add x3, x1, x2 => 34+55=89
    RAM[41] = 32'h003026A3; // sw x3, 44(x0) => 89
    RAM[42] = 32'h002000B3; // add x1, x0, x2 => x1=55
    RAM[43] = 32'h00300133; // add x2, x0, x3 => x2=89

    RAM[44] = 32'h002081B3; // add x3, x1, x2 => 55+89=144
    RAM[45] = 32'h003028A3; // sw x3, 48(x0) => 144
    RAM[46] = 32'h002000B3; // add x1, x0, x2 => x1=89
    RAM[47] = 32'h00300133; // add x2, x0, x3 => x2=144

    RAM[48] = 32'h002081B3; // add x3, x1, x2 => 89+144=233
    RAM[49] = 32'h00302AA3; // sw x3, 52(x0) => 233
    RAM[50] = 32'h002000B3; // add x1, x0, x2 => x1=144
    RAM[51] = 32'h00300133; // add x2, x0, x3 => x2=233

    RAM[52] = 32'h002081B3; // add x3, x1, x2 => 144+233=377
    RAM[53] = 32'h00302CA3; // sw x3, 56(x0) => 377
    RAM[54] = 32'h002000B3; // add x1, x0, x2 => x1=233
    RAM[55] = 32'h00300133; // add x2, x0, x3 => x2=377

    RAM[56] = 32'h002081B3; // add x3, x1, x2 => 233+377=610
    RAM[57] = 32'h00302EA3; // sw x3, 60(x0) => 610
    RAM[58] = 32'h002000B3; // add x1, x0, x2 => x1=377
    RAM[59] = 32'h00300133; // add x2, x0, x3 => x2=610

    RAM[60] = 32'h002081B3; // add x3, x1, x2 => 377+610=987
    RAM[61] = 32'h00302023; // sw x3, 64(x0) => 987
    RAM[62] = 32'h002000B3; // add x1, x0, x2 => x1=610
    RAM[63] = 32'h00300133; // add x2, x0, x3 => x2=987

    RAM[64] = 32'h002081B3; // add x3, x1, x2 => 610+987=1597
    RAM[65] = 32'h00302223; // sw x3, 68(x0) => 1597
    RAM[66] = 32'h002000B3; // add x1, x0, x2 => x1=987
    RAM[67] = 32'h00300133; // add x2, x0, x3 => x2=1597

    RAM[68] = 32'h002081B3; // add x3, x1, x2 => 987+1597=2584
    RAM[69] = 32'h00302423; // sw x3, 72(x0) => 2584
    RAM[70] = 32'h002000B3; // add x1, x0, x2 => x1=1597
    RAM[71] = 32'h00300133; // add x2, x0, x3 => x2=2584

    RAM[72] = 32'h002081B3; // add x3, x1, x2 => 1597+2584=4181
    RAM[73] = 32'h00302623; // sw x3, 76(x0) => 4181
    RAM[74] = 32'h002000B3; // add x1, x0, x2 => x1=2584
    RAM[75] = 32'h00300133; // add x2, x0, x3 => x2=4181
    
    RAM[76] = 32'h002081B3; // add x3, x1, x2 => 2584+4181=6765
    RAM[77] = 32'h00302423; // sw x3, 80(x0) => 6765
    RAM[78] = 32'h00000093; // addi x1, x0, 0
    RAM[79] = 32'h00100113; // addi x2, x0, 1
    RAM[80] = 32'hEC1FF0EF; // jal x0, -320 (go back to RAM[0])
   
    end
endmodule