module controlpath();

endmodule