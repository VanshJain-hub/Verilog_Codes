module mux_using2to1(
    input a,b,c,d
);